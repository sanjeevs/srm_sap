//
// Package for blockA backdoor logic.
//

package blockA_backdoor_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import srm_pkg::*;
  `include "blockA_backdoor_adapter.svh"
  `include "blockA_backdoor_handle.svh"
endpackage

