//
// Package for the pio agent
//

package pio_agent_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import srm_pkg::*;
  `include "pio_xact.svh"
  `include "pio_seq_lib.svh"
  `include "pio_driver.svh"
  `include "pio_sequencer.svh"
  `include "pio_agent_config.svh"
  `include "pio_bus_adapter.svh"
  `include "pio_bus_handle.svh"
  `include "pio_agent.svh"
endpackage

