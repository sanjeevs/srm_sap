//
// Package for sap1 register model
//
package sap1_srm_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import srm_pkg::*;
  import sap1_srm_model_pkg::*;

  `include "srm_frontdoor_handle.svh"
  `include "sap1_srm_reg_sequence.svh"
endpackage
