//
// Package for sap2_srm_model
//
`ifndef INCLUDED_sap2_srm_model_pkg
`define INCLUDED_sap2_srm_model_pkg

package sap2_srm_model_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import srm_pkg::*;

  import blockA_srm_model_pkg::*;
  import sap1_srm_model_pkg::*;
  `include "sap2_srm_model.svh"
endpackage

`endif
