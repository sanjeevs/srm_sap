//
// Package for blockA_srm_constr_model
//
`ifndef INCLUDED_blockA_srm_constr_pkg
`define INCLUDED_blockA_srm_constr_pkg

package blockA_srm_constr_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import srm_pkg::*;
  import blockA_srm_model_pkg::*;

  `include "blockA_srm_constr.svh"
endpackage

`endif
