//
// Package for the host agent
//

package host_agent_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "host_xact.svh"
  `include "host_seq_lib.svh"
  `include "host_driver.svh"
  `include "host_sequencer.svh"
  `include "host_agent.svh"
endpackage

