//
// Package for the sap2 env
//

package sap2_env_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import srm_pkg::*; 
  import host_agent_pkg::*;
  import pio_agent_pkg::*;
  `include "sap2_env_config.svh"
  `include "sap2_env.svh"
endpackage
