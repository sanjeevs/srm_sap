//
// Package for the blockA reg sequences.
//

package blockA_srm_reg_sequences_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import srm_pkg::*; 
  import blockA_srm_model_pkg::*;   
  `include "blockA_srm_reg_sequence.svh"
  `include "blockA_srm_table_sequence.svh"
endpackage
