//
// Package for sap1_srm_model
//
`ifndef INCLUDED_sap1_srm_model_pkg
`define INCLUDED_sap1_srm_model_pkg

package sap1_srm_model_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import srm_pkg::*;

  `include "sap1_srm_model.svh"
endpackage

`endif
