//
// Package for blockA_srm_model
//
`ifndef INCLUDED_blockA_srm_model_pkg
`define INCLUDED_blockA_srm_model_pkg

package blockA_srm_model_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import srm_pkg::*;

  `include "blockA_srm_model.svh"
endpackage

`endif
