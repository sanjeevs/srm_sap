//
// Package for the host agent
//

package host_agent_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import srm_pkg::*;
  `include "host_xact.svh"
  `include "host_seq_lib.svh"
  `include "host_driver.svh"
  `include "host_sequencer.svh"
  `include "host_agent_config.svh"
  `include "host_agent.svh"
  `include "host_bus_adapter.svh"
endpackage

